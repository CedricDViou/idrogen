library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_arith.all;
use IEEE.STD_LOGIC_unsigned.all;
use work.pack_ipv4_types.all;
use work.ipbus.all;

--library unisim;
--use unisim.VComponents.all;

entity ipbus_1G is
    generic (
        IN_SIMULATION        : BOOLEAN                       := false;
        SIMUL_DST_MAC_NUMBER : STD_LOGIC_VECTOR(47 downto 0) := x"AAAA_BBBB_CCCC";
        CLOCK_FREQ           : INTEGER                       := 125000000; -- freq of data_in_clk -- needed to timout cntr
        DHCP_CLOCK_FREQ      : INTEGER                       := 125000000; -- freq of data_in_clk -- needed to timout cntr
        LEASE_TIME_TO_REQ    : INTEGER                       := 60;        -- lease time request (in sec)
        ARP_TIMEOUT          : INTEGER                       := 60;        -- ARP response timeout (s)
        ARP_MAX_PKT_TMO      : INTEGER                       := 5;         -- # wrong nwk pkts received before set error
        MAX_ARP_ENTRIES      : INTEGER                       := 255        -- max entries in the ARP store
    );
    port (
        clk125                          : in  STD_LOGIC;
        rst_125                         : in  STD_LOGIC;
        phy_rstb                        : out STD_LOGIC;
        rx_gbt                          : in  STD_LOGIC;
        tx_gbt                          : out STD_LOGIC;
        spi_interface_address           : in  STD_LOGIC_VECTOR(26 downto 0);  -- address
        spi_interface_byte_enable       : in  STD_LOGIC_VECTOR(3 downto 0);   -- byte_enable
        spi_interface_read              : in  STD_LOGIC;                      -- read
        spi_interface_write             : in  STD_LOGIC;                      -- write
        spi_interface_write_data        : in  STD_LOGIC_VECTOR(31 downto 0);  -- write_data
        spi_interface_acknowledge       : out STD_LOGIC;                      -- acknowledge
        spi_interface_read_data         : out STD_LOGIC_VECTOR(31 downto 0);  -- read_data
        uc_interrupt                    : out STD_LOGIC;
        ipbus_uart_rxd                  : in  STD_LOGIC;                      -- uart.rxd
        ipbus_uart_txd                  : out STD_LOGIC                       --     .txd
    );
end ipbus_1G;

architecture RTL of ipbus_1G is

    constant nb_src : NATURAL := 2;
    component UDP_Complete
        generic (
            IN_SIMULATION        : BOOLEAN                       := false;
            SIMUL_DST_MAC_NUMBER : STD_LOGIC_VECTOR(47 downto 0) := x"AAAA_BBBB_CCCC";
            CLOCK_FREQ           : INTEGER                       := 125000000; -- freq of data_in_clk -- needed to timout cntr
            ARP_TIMEOUT          : INTEGER                       := 60;        -- ARP response timeout (s)
            ARP_MAX_PKT_TMO      : INTEGER                       := 5;         -- # wrong nwk pkts received before set error
            MAX_ARP_ENTRIES      : INTEGER                       := 255        -- max entries in the ARP store
        );
        port (
            -- UDP TX signals
            udp_tx_start          : in STD_LOGIC;   -- indicates req to tx UDP
            udp_txi               : in udp_tx_type; -- UDP tx cxns
            udp_tx_result         : out STD_LOGIC_VECTOR (1 downto 0);-- tx status (changes during transmission)
            udp_tx_data_out_ready : out STD_LOGIC; -- indicates udp_tx is ready to take data

            -- UDP RX signals
            udp_rx_start : out STD_LOGIC; -- indicates receipt of udp header
            udp_rxo      : out udp_rx_type;

            -- IP RX signals
            ip_rx_hdr : out ipv4_rx_header_type;

            -- system signals
            clk125          : in STD_LOGIC;
            reset           : in STD_LOGIC;
            our_ip_address  : in STD_LOGIC_VECTOR (31 downto 0);
            our_mac_address : in STD_LOGIC_VECTOR (47 downto 0);
            gateway         : in STD_LOGIC_VECTOR(31 downto 0);
            netmask         : in STD_LOGIC_VECTOR(31 downto 0);
            control         : in udp_control_type;

            -- status signals
            arp_pkt_count : out STD_LOGIC_VECTOR(7 downto 0); -- count of arp pkts received
            ip_pkt_count  : out STD_LOGIC_VECTOR(7 downto 0); -- number of IP pkts received for us

            -- gmii TX interface
            --     gmii_gtx_clk : out STD_LOGIC; -- must be generated with appropriate system
            gmii_tx_en : out STD_LOGIC;
            gmii_tx_er : out STD_LOGIC;
            gmii_txd   : out STD_LOGIC_VECTOR(7 downto 0);

            -- gmii RX interface
            gmii_rx_clk : in STD_LOGIC;
            gmii_rx_dv  : in STD_LOGIC;
            gmii_rx_er  : in STD_LOGIC;
            gmii_rxd    : in STD_LOGIC_VECTOR(7 downto 0)
        );
    end component;

    component dhcp_client
        generic (
            CLOCK_FREQ        : INTEGER := 125000000; -- freq of data_in_clk -- needed to timout cntr
            LEASE_TIME_TO_REQ : INTEGER := 3600       -- lease time request (in sec)
        );
        port (
            -- system signals
            clk             : in STD_LOGIC;
            reset           : in STD_LOGIC;
            our_mac_address : in STD_LOGIC_VECTOR (47 downto 0);

            -- UDP TX signals
            udp_tx_start          : out STD_LOGIC;                    -- indicates req to tx UDP
            udp_txi               : out udp_tx_type;                  -- UDP tx cxns
            udp_tx_result         : in STD_LOGIC_VECTOR (1 downto 0); -- tx status (changes during transmission)
            udp_tx_data_out_ready : in STD_LOGIC;                     -- indicates udp_tx is ready to take data

            -- UDP RX signals
            udp_rx_start : in STD_LOGIC; -- indicates receipt of udp header
            udp_rxo      : in udp_rx_type;

            gateway              : out STD_LOGIC_VECTOR(31 downto 0);
            netmask              : out STD_LOGIC_VECTOR(31 downto 0);
            allocated_ip_address : out STD_LOGIC_VECTOR (31 downto 0)

        );
    end component;

    component ipbus_qsys is
        port (
            clk_clk                                                 : in  STD_LOGIC                      := 'X';              -- clk
            ipbus_avallon_master_1_ipbread_ipbus_read_readdata      : out STD_LOGIC_VECTOR(31 downto 0)  := (others => 'X');  -- ipbus_read_readdata
            ipbus_avallon_master_1_ipbread_ipbus_read_ack           : out STD_LOGIC                      := 'X';              -- ipbus_read_ack
            ipbus_avallon_master_1_ipbread_ipbus_read_err           : out STD_LOGIC                      := 'X';              -- ipbus_read_err
            ipbus_avallon_master_1_ipbuswrite_ipbus_write_addr      : in  STD_LOGIC_VECTOR(31 downto 0)  := (others => 'X');  -- ipbus_write_addr
            ipbus_avallon_master_1_ipbuswrite_ipbus_write_writedata : in  STD_LOGIC_VECTOR(31 downto 0)  := (others => 'X');  -- ipbus_write_writedata
            ipbus_avallon_master_1_ipbuswrite_ipbus_write_strobe    : in  STD_LOGIC                      := 'X';              -- ipbus_write_strobe
            ipbus_avallon_master_1_ipbuswrite_ipbus_write_write     : in  STD_LOGIC                      := 'X';              -- ipbus_write_write
            reset_reset                                             : in  STD_LOGIC                      := 'X';              -- reset
            spi_interface_address                                   : in  STD_LOGIC_VECTOR(26 downto 0)  := (others => 'X');
            spi_interface_byte_enable                               : in  STD_LOGIC_VECTOR(3 downto 0)   := (others => 'X');
            spi_interface_read                                      : in  STD_LOGIC                      := 'X';
            spi_interface_write                                     : in  STD_LOGIC                      := 'X';
            spi_interface_write_data                                : in  STD_LOGIC_VECTOR(31 downto 0)  := (others => 'X');
            spi_interface_acknowledge                               : out STD_LOGIC;
            spi_interface_read_data                                 : out STD_LOGIC_VECTOR(31 downto 0);
            ipbus_to_uart_rxd                                       : in  STD_LOGIC                     := 'X';               -- uart.rxd
            ipbus_to_uart_txd                                       : out STD_LOGIC;                                          --     .txd
            spi_export                                              : out STD_LOGIC_VECTOR(7 downto 0);                       -- export
            mac_address_export                                      : out STD_LOGIC_VECTOR(7 downto 0);
            bridge_uart_address                                     : in  STD_LOGIC_VECTOR(5 downto 0)  := (others => 'X'); -- address
            bridge_uart_byte_enable                                 : in  STD_LOGIC_VECTOR(3 downto 0)  := (others => 'X'); -- byte_enable
            bridge_uart_read                                        : in  STD_LOGIC                     := 'X';             -- read
            bridge_uart_write                                       : in  STD_LOGIC                     := 'X';             -- write
            bridge_uart_write_data                                  : in  STD_LOGIC_VECTOR(31 downto 0) := (others => 'X'); -- write_data
            bridge_uart_acknowledge                                 : out STD_LOGIC;                                        -- acknowledge
            bridge_uart_read_data                                   : out STD_LOGIC_VECTOR(31 downto 0)                     -- read_data
        );
    end component ipbus_qsys;

    component wr_monitor
        port (
            clock                   : in  STD_LOGIC;
            nreset                  : in  STD_LOGIC;
            bridge_uart_acknowledge : in  STD_LOGIC;
            bridge_uart_read_data   : in  STD_LOGIC_VECTOR (31 downto 0);
            bridge_uart_read        : out STD_LOGIC;
            bridge_uart_write       : out STD_LOGIC;
            bridge_uart_byte_enable : out STD_LOGIC_VECTOR ( 3 downto 0);
            bridge_uart_address     : out STD_LOGIC_VECTOR ( 5 downto 0);
            bridge_uart_write_data  : out STD_LOGIC_VECTOR (31 downto 0)
        );
    end component;


    component MyGbt
        port (
            pll_refclk        : in  STD_LOGIC;
            reset             : in  STD_LOGIC;
            rx_ready          : out STD_LOGIC;
            tx_ready          : out STD_LOGIC;
            rx_gbt            : in  STD_LOGIC;
            tx_gbt            : out STD_LOGIC;
            rx_is_lockedtoref : out STD_LOGIC;
            rx_parallel_data  : out STD_LOGIC_VECTOR(7 downto 0);
            tx_parallel_data  : in  STD_LOGIC_VECTOR(7 downto 0);
            rx_datak          : out STD_LOGIC;
            tx_datak          : in  STD_LOGIC;
            rx_errdetect      : out STD_LOGIC;
            rx_disperr        : out STD_LOGIC;
            rx_runningdisp    : out STD_LOGIC;
            rx_patterndetect  : out STD_LOGIC;
            rx_rmfifostatus   : out STD_LOGIC_VECTOR(1 downto 0);
            rx_syncstatus     : out STD_LOGIC;
            tx_clk            : out STD_LOGIC;
            rx_clk            : out STD_LOGIC
        );
    end component;

    component ipbus_main
        generic (
            -- Number of RX and TX buffers is 2**BUFWIDTH
            BUFWIDTH : NATURAL := 4;
            -- Number of address bits within each buffer in UDP I/F
            -- Size of each buffer is 2**ADDRWIDTH --MAXIMUM is 14 bit
            ADDRWIDTH : NATURAL := 9;
            -- UDP port for IPbus traffic in this instance of UDP I/F
            IPBUSPORT : STD_LOGIC_VECTOR(15 downto 0) := x"C351"
        );
        port (
            mac_clk    : in STD_LOGIC; -- Ethernet MAC clock (125MHz)
            rst_macclk : in STD_LOGIC; -- MAC clock domain sync reset

            -- UDP RX signals
            udp_rx_start : in STD_LOGIC; -- indicates receipt of udp header
            udp_rxo      : in udp_rx_type;

            -- UDP TX signals
            udp_tx_start          : out STD_LOGIC;                    -- indicates req to tx UDP
            udp_txi               : out udp_tx_type;                  -- UDP tx cxns
            udp_tx_result         : in STD_LOGIC_VECTOR (1 downto 0); -- tx status (changes during transmission)
            udp_tx_data_out_ready : in STD_LOGIC;                     -- indicates udp_tx is ready to take data

            -- ipb interface
            ipb_clk : in STD_LOGIC; -- IPbus clock
            rst_ipb : in STD_LOGIC; -- IPbus clock domain sync reset
            ipb_out : out ipb_wbus;
            ipb_in  : in ipb_rbus
        );
    end component;

    component udp_tx_arbitrer
        generic (
            nb_src : NATURAL
        );
        port (
            mac_clk    : in STD_LOGIC; -- Ethernet MAC clock (125MHz)
            rst_macclk : in STD_LOGIC; -- MAC clock domain sync reset

            -- UDP result TX signals
            src_udp_tx_start          : in STD_LOGIC_VECTOR(0 to nb_src - 1);
            src_udp_tx                : in udp_tx_vect_type(0 to nb_src - 1);
            src_udp_tx_result         : out Array2bit_ip(0 to nb_src - 1);     -- tx status (changes during transmission)
            src_udp_tx_data_out_ready : out STD_LOGIC_VECTOR(0 to nb_src - 1); -- indicates udp_tx is ready to take data

            -- UDP result TX signals
            arb_udp_tx_start          : out STD_LOGIC; -- indicates req to tx UDP
            arb_udp_txi               : out udp_tx_type;
            arb_udp_tx_result         : in STD_LOGIC_VECTOR (1 downto 0); -- tx status (changes during transmission)
            arb_udp_tx_data_out_ready : in STD_LOGIC                      -- indicates udp_tx is ready to take data
        );
    end component udp_tx_arbitrer;

    --UDP/IPBUS interconnection
    signal udp_tx_start_ipbus          : STD_LOGIC; -- indicates req to tx UDP
    signal udp_txi_ipbus               : udp_tx_type;
    signal udp_tx_result_ipbus         : STD_LOGIC_VECTOR (1 downto 0);-- tx status (changes during transmission)
    signal udp_tx_data_out_ready_ipbus : STD_LOGIC; -- indicates udp_tx is ready to take data

    signal udp_rx_start : STD_LOGIC; -- indicates receipt of udp header
    signal udp_rxo      : udp_rx_type;

    signal control : udp_control_type;

    signal rx_clk, rx_clk_io : STD_LOGIC;
    signal txd_e, rxd_r      : STD_LOGIC_VECTOR(7 downto 0);
    signal tx_en_e, tx_er_e  : STD_LOGIC;
    signal rx_dv_r, rx_er_r  : STD_LOGIC;
    signal gmii_rxd_del      : STD_LOGIC_VECTOR(7 downto 0);
    signal gmii_rx_dv_del    : STD_LOGIC;
    signal gmii_rx_er_del    : STD_LOGIC;
    signal our_ip_address    : STD_LOGIC_VECTOR (31 downto 0);
    signal our_mac_address   : STD_LOGIC_VECTOR (47 downto 0);

    -- IPBUS connection
    signal ipb_out     : ipb_wbus;
    signal ipb_in      : ipb_rbus;
    signal gmii_rx_clk : STD_LOGIC;
    signal gateway     : STD_LOGIC_VECTOR(31 downto 0);
    signal netmask     : STD_LOGIC_VECTOR(31 downto 0);

    -- gmii TX interface
    signal gmii_tx_en : STD_LOGIC;
    signal gmii_tx_er : STD_LOGIC;
    signal gmii_txd   : STD_LOGIC_VECTOR(7 downto 0);

    -- gmii RX interface
    signal gmii_rx_dv : STD_LOGIC;

    signal udp_tx_start_dhcp          : STD_LOGIC;
    signal udp_txi_dhcp               : udp_tx_type;
    signal udp_tx_result_dhcp         : STD_LOGIC_VECTOR (1 downto 0);
    signal udp_tx_data_out_ready_dhcp : STD_LOGIC;

    signal udp_tx_start_arb          : STD_LOGIC;
    signal udp_txi_arb               : udp_tx_type;
    signal udp_tx_result_arb         : STD_LOGIC_VECTOR (1 downto 0);
    signal udp_tx_data_out_ready_arb : STD_LOGIC;

    signal src_udp_tx_start          : STD_LOGIC_VECTOR(0 to nb_src - 1);
    signal src_udp_tx                : udp_tx_vect_type(0 to nb_src - 1);
    signal src_udp_tx_result         : Array2bit_ip(0 to nb_src - 1);     -- tx status (changes during transmission)
    signal src_udp_tx_data_out_ready : STD_LOGIC_VECTOR(0 to nb_src - 1); -- indicates udp_tx is ready to take data

    signal spi_export                : STD_LOGIC_VECTOR (7 downto 0);
    signal mac_address_export        : STD_LOGIC_VECTOR (7 downto 0);

    signal bridge_uart_read          : STD_LOGIC;
    signal bridge_uart_write         : STD_LOGIC;
    signal bridge_uart_acknowledge   : STD_LOGIC;
    signal bridge_uart_byte_enable   : STD_LOGIC_VECTOR ( 3 downto 0);
    signal bridge_uart_address       : STD_LOGIC_VECTOR ( 5 downto 0);
    signal bridge_uart_read_data     : STD_LOGIC_VECTOR (31 downto 0);
    signal bridge_uart_write_data    : STD_LOGIC_VECTOR (31 downto 0);
    
begin

    -------------------------------------------------------------------------------
    -- UDP connection
    -------------------------------------------------------------------------------
    lbl_UDP : UDP_Complete generic map(
        IN_SIMULATION        => IN_SIMULATION,
        SIMUL_DST_MAC_NUMBER => SIMUL_DST_MAC_NUMBER,

        CLOCK_FREQ      => CLOCK_FREQ,
        ARP_TIMEOUT     => ARP_TIMEOUT,
        ARP_MAX_PKT_TMO => ARP_MAX_PKT_TMO,
        MAX_ARP_ENTRIES => MAX_ARP_ENTRIES
    )
    port map(
        -- UDP TX signals
        udp_tx_start          => udp_tx_start_arb,          -- udp_tx_start,
        udp_txi               => udp_txi_arb,               -- udp_txi,
        udp_tx_result         => udp_tx_result_arb,         -- udp_tx_result,
        udp_tx_data_out_ready => udp_tx_data_out_ready_arb, -- udp_tx_data_out_ready,

        -- UDP RX signals
        udp_rx_start => udp_rx_start,
        udp_rxo      => udp_rxo,

        -- IP RX signals
        ip_rx_hdr => open,

        -- system signals
        clk125          => clk125,
        reset           => rst_125,
        our_ip_address  => our_ip_address,
        our_mac_address => our_mac_address,
        gateway         => gateway,
        netmask         => netmask,
        control         => control,

        -- status signals
        arp_pkt_count => open,
        ip_pkt_count  => open,

        -- gmii TX interface
        -- gmii_gtx_clk : out STD_LOGIC; -- must be generated with appropriate system
        gmii_txd   => txd_e,
        gmii_tx_en => tx_en_e,
        gmii_tx_er => tx_er_e,

        -- gmii RX interface
        gmii_rx_clk => rx_clk,
        gmii_rxd    => rxd_r,
        gmii_rx_dv  => rx_dv_r,
        gmii_rx_er  => '0');

    our_mac_address                              <= x"00228f5555" & mac_address_export;
    control.ip_controls.arp_controls.clear_cache <= '0';

    -------------------------------------------------------------------------------
    --  dhcp block
    -------------------------------------------------------------------------------
    lbl_dhcp : dhcp_client generic map(
        CLOCK_FREQ        => DHCP_CLOCK_FREQ,
        LEASE_TIME_TO_REQ => LEASE_TIME_TO_REQ
    )
    port map(
        -- system signals
        clk             => clk125,
        reset           => rst_125,
        our_mac_address => our_mac_address,

        -- UDP TX signals
        udp_tx_start          => udp_tx_start_dhcp,          --udp_tx_start,
        udp_txi               => udp_txi_dhcp,               --udp_txi,
        udp_tx_result         => udp_tx_result_dhcp,         --udp_tx_result,
        udp_tx_data_out_ready => udp_tx_data_out_ready_dhcp, --udp_tx_data_out_ready,

        -- UDP RX signals
        udp_rx_start => udp_rx_start,
        udp_rxo      => udp_rxo,

        gateway              => gateway,
        netmask              => netmask,
        allocated_ip_address => our_ip_address
    );

    -------------------------------------------------------------------------------
    -- IPBUS block
    -------------------------------------------------------------------------------
    lbl_ipbus : ipbus_main generic map(
        -- Number of RX and TX buffers is 2**BUFWIDTH
        BUFWIDTH => 4,
        -- Number of address bits within each buffer in UDP I/F
        -- Size of each buffer is 2**ADDRWIDTH --MAXIMUM is 14 bit
        ADDRWIDTH => 9,
        -- UDP port for IPbus traffic in this instance of UDP I/F
        IPBUSPORT => x"C351"
    )
    port map(
        mac_clk    => clk125,
        rst_macclk => rst_125,

        -- UDP RX signals
        udp_rx_start => udp_rx_start,
        udp_rxo      => udp_rxo,

        -- UDP TX signals
        udp_tx_start          => udp_tx_start_ipbus,
        udp_txi               => udp_txi_ipbus,
        udp_tx_result         => udp_tx_result_ipbus,
        udp_tx_data_out_ready => udp_tx_data_out_ready_ipbus,

        -- ipb interface
        ipb_clk => clk125,
        rst_ipb => rst_125,
        ipb_out => ipb_out,
        ipb_in  => ipb_in
    );

    -------------------------------------------------------------------------------
    -- IPBUS/UDP arbitrer
    -------------------------------------------------------------------------------
    lbl_udp_arb : udp_tx_arbitrer generic map(nb_src)
    port map(
        mac_clk    => clk125,
        rst_macclk => rst_125,

        src_udp_tx_start          => src_udp_tx_start,
        src_udp_tx                => src_udp_tx,
        src_udp_tx_result         => src_udp_tx_result,
        src_udp_tx_data_out_ready => src_udp_tx_data_out_ready,

        -- UDP result TX signals
        arb_udp_tx_start          => udp_tx_start_arb,
        arb_udp_txi               => udp_txi_arb,
        arb_udp_tx_result         => udp_tx_result_arb,
        arb_udp_tx_data_out_ready => udp_tx_data_out_ready_arb
    );

    -- UDP result TX signals (ipbus)
    src_udp_tx_start(0)         <= udp_tx_start_ipbus;
    src_udp_tx(0)               <= udp_txi_ipbus;
    udp_tx_result_ipbus         <= src_udp_tx_result(0);
    udp_tx_data_out_ready_ipbus <= src_udp_tx_data_out_ready(0);

    -- UDP result TX signals (dhcp)
    src_udp_tx_start(1)        <= udp_tx_start_dhcp;
    src_udp_tx(1)              <= udp_txi_dhcp;
    udp_tx_result_dhcp         <= src_udp_tx_result(1);
    udp_tx_data_out_ready_dhcp <= src_udp_tx_data_out_ready(1);

    u0 : component ipbus_qsys
        port map(
            clk_clk                                                 => clk125,             --                               clk.clk
            ipbus_avallon_master_1_ipbread_ipbus_read_readdata      => ipb_in.ipb_rdata,   --    ipbus_avallon_master_0_ipbread.ipbus_read_readdata
            ipbus_avallon_master_1_ipbread_ipbus_read_ack           => ipb_in.ipb_ack,     --                                  .ipbus_read_ack
            ipbus_avallon_master_1_ipbread_ipbus_read_err           => ipb_in.ipb_err,     --                                  .ipbus_read_err
            ipbus_avallon_master_1_ipbuswrite_ipbus_write_addr      => ipb_out.ipb_addr,   -- ipbus_avallon_master_0_ipbuswrite.ipbus_write_addr
            ipbus_avallon_master_1_ipbuswrite_ipbus_write_writedata => ipb_out.ipb_wdata,  --                                  .ipbus_write_writedata
            ipbus_avallon_master_1_ipbuswrite_ipbus_write_strobe    => ipb_out.ipb_strobe, --                                  .ipbus_write_strobe
            ipbus_avallon_master_1_ipbuswrite_ipbus_write_write     => ipb_out.ipb_write,  --                                  .ipbus_write_write
            reset_reset                                             => rst_125,            --                             reset.reset
            spi_interface_address                                   => spi_interface_address,
            spi_interface_byte_enable                               => spi_interface_byte_enable,
            spi_interface_read                                      => spi_interface_read,
            spi_interface_write                                     => spi_interface_write,
            spi_interface_write_data                                => spi_interface_write_data,
            spi_interface_acknowledge                               => spi_interface_acknowledge,
            spi_interface_read_data                                 => spi_interface_read_data,
            ipbus_to_uart_rxd                                       => ipbus_uart_rxd,
            ipbus_to_uart_txd                                       => ipbus_uart_txd,
            spi_export                                              => spi_export,       --         pio_0_external_connection.export
            mac_address_export                                      => mac_address_export,
            bridge_uart_address                                     => bridge_uart_address,
            bridge_uart_byte_enable                                 => bridge_uart_byte_enable,
            bridge_uart_read                                        => bridge_uart_read,
            bridge_uart_write                                       => bridge_uart_write,
            bridge_uart_write_data                                  => bridge_uart_write_data,
            bridge_uart_acknowledge                                 => bridge_uart_acknowledge,
            bridge_uart_read_data                                   => bridge_uart_read_data
        );

    wr_monitor_inst : wr_monitor
        port map (
            clock                   => clk125,
            nreset                  => rst_125,
            bridge_uart_acknowledge => bridge_uart_acknowledge,
            bridge_uart_read_data   => bridge_uart_read_data,
            bridge_uart_read        => bridge_uart_read,
            bridge_uart_write       => bridge_uart_write,
            bridge_uart_byte_enable => bridge_uart_byte_enable,
            bridge_uart_address     => bridge_uart_address,
            bridge_uart_write_data  => bridge_uart_write_data
        );

    uc_interrupt <= spi_export(0);

    -------------------------------------------------------------------------------
    -- IO interface
    -------------------------------------------------------------------------------
    phy_rstb <= '1';

    rx_clk_io <= gmii_rx_clk;
    rx_clk    <= gmii_rx_clk;
    process (rx_clk_io) -- FFs for incoming GMII data (need to be IOB FFs)
    begin
        if rising_edge(rx_clk_io) then
            rxd_r   <= gmii_rxd_del;
            rx_dv_r <= gmii_rx_dv_del;
            rx_er_r <= gmii_rx_er_del; -- Que faire de ce signal?
        end if;
    end process;

    process (clk125) -- FFs for outgoing GMII data (need to be IOB FFs)
    begin
        if rising_edge(clk125) then
            gmii_txd   <= txd_e;
            gmii_tx_en <= tx_en_e;
            gmii_tx_er <= tx_er_e; --Que faire avec ce signal ?
        end if;
    end process;

    -------------------------------------------------------------------------------
    -- Internal Phy interface
    -------------------------------------------------------------------------------
    mygbt_inst : mygbt
    port map(
        pll_refclk        => clk125,
        reset             => rst_125,
        rx_ready          => open,
        tx_ready          => open,
        rx_gbt            => rx_gbt,
        tx_gbt            => tx_gbt,
        rx_is_lockedtoref => open,
        rx_parallel_data  => gmii_rxd_del,
        tx_parallel_data  => gmii_txd,
        rx_datak          => gmii_rx_dv_del,
        tx_datak          => gmii_tx_en,
        rx_errdetect      => open,
        rx_disperr        => open,
        rx_runningdisp    => open,
        rx_patterndetect  => open,
        rx_rmfifostatus   => open,
        rx_syncstatus     => open,
        tx_clk            => open,
        rx_clk            => gmii_rx_clk
    );

end RTL;