// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.1.0 Build 222 09/21/2018 SJ Pro Edition
// Created on Fri Feb 18 19:44:24 2022

// synthesis message_off 10175

//`timescale 1ns/1ns

//! State Machine interface between SPI slave module and Avallon External Bus

module SPI_SM (
    nreset, clock, ack, bit_cnt[6:0], csn, read_data_from_avallon[31:0], data_from_spi[31:0],
    address[31:0], read, write, byte_enable[3:0], read_data_to_spi[31:0], write_data_to_avallon[31:0]);

    input 			nreset;                 //! Reset actif a l'etat bas
    input 			clock;                  //! Horloge
    input 			ack;                    //! Signal d'acknoledge provenant du bus avalon pour signaler que l'operation de lecture/ecriture est terminee.
    input 			csn;                    //! Chip select
    //input 			rw;                 // Bit de lecture/ecriture
	input  [6:0] 	bit_cnt;                //! Position dans la trame SPI
    input [31:0] 	read_data_from_avallon; //! Donnee recue du bus avallon
    input [31:0] 	data_from_spi;    		//! Donnee recue du bus SPI
	
    tri0 		nreset;
    tri0 		ack;
    tri0 		csn;
//    tri0 		rw;
	tri0  [6:0] bit_cnt;
    tri0 [31:0] read_data_from_avallon;
    tri0 [31:0] data_from_spi;
	
    output reg 			read;                   //! Signal positionne a "1" pour indiquer au bus avallon que l'on souhaite realiser une operation de lecture
    output reg			write;                  //! Signal positionne a "1" pour indiquer au bus avallon que l'on souhaite realiser une operation d'ecriture
    output reg  [3:0] 	byte_enable;            //! Indique les octets a lire/ecrire dans le mot de 32 bits
    output reg [31:0] 	read_data_to_spi;       //! Donnee de lecture a transmettre au processus SPI
    output reg [31:0] 	write_data_to_avallon;  //! Donnee d'ecriture a transmettre a l'interface avallon
	output reg [31:0] 	address;				//! Adresse de lecture/ecriture sur le bus avallon
	
	reg  [6:0] 	reg_fstate; //! Registre d'etat
    
    reg 		ack_synchro;                    
	reg  [6:0] 	bit_cnt_synchro;                //! Resynchronisation du registre bit_cnt
    reg [31:0] 	data_from_spi_synchro;    		//! Resynchronisation du registre data_from_spi
    reg [31:0] 	read_data_from_avallon_synchro; //! Resynchronisation du registre read_data_from_avallon

    //! Resynchronisation des signaux d'entrée sur le nouveau domaine d'horloge
    always @(posedge clock or negedge nreset or posedge csn)
    begin : sync_prosses
        if (~nreset || csn) begin
            ack_synchro 					<=  1'b0;
            bit_cnt_synchro      		    <=  7'd0;
			data_from_spi_synchro 		    <= 32'h0;
            read_data_from_avallon_synchro 	<= 32'h0;
        end
        else begin
            ack_synchro 					<= ack;
            bit_cnt_synchro      		    <= bit_cnt;
			data_from_spi_synchro 		    <= data_from_spi;
            read_data_from_avallon_synchro 	<= read_data_from_avallon;
        end
    end
	
	// IDLE 				= 7'd0
	// GET ADDRESS 			= 7'd1
	// READ_AVALON 			= 7'd2
	// SEND_SPI				= 7'd4
	// GET_SPI				= 7'd8
	// WRITE_AVALON 		= 7'd16
	// WAIT_WRITE_END_FRAME = 7'd32
	// WAIT_READ_END_FRAME 	= 7'd64
	
    //! State Machine process : update state
    //! fsm_extract
	always @(posedge clock or negedge nreset or posedge csn)
    begin : state_machine_interface
        if (~nreset || csn) begin
            reg_fstate [6:0]		<=  7'd0;
            read 					<=  1'b0;
            write 					<=  1'b0;
            byte_enable 			<=  4'h0;
            address 				<= 32'h0;
			read_data_to_spi 		<= 32'h0;
            write_data_to_avallon 	<= 32'h0;
        end
        else begin
            case (reg_fstate)
                7'd0: begin
					reg_fstate [6:0]		<=  7'd1;   // Sortie de l'etat IDLE et debut de la lecture de l'adresse
					read 					<=  1'b0;
					write 					<=  1'b0;
					byte_enable 			<=  4'h0;
					address 				<= 32'h0;
					read_data_to_spi 		<= 32'h0;
					write_data_to_avallon 	<= 32'h0;
                end
                7'd1: begin	
                    if (bit_cnt_synchro==7'h20) begin
                        address [31:0]	<= {1'b0, data_from_spi_synchro[30:0]};
                        if (data_from_spi_synchro[31])
                            reg_fstate [6:0] 	<= 7'd2;    // L'adresse est recue et on commence la lecture du bus avallon
                        else
                            reg_fstate [6:0] 	<= 7'd8;    // L'adresse est recue et on commence la reception de la donnee a ecrire
                    end
                    else begin
                        reg_fstate [6:0] 	<= 7'd1;
                        address             <= address; 
					end
                end
                7'd2: begin
                    // Operation de lecture : les registres "read" et "byte_enable" sont actif pour lancer la lecture au niveau du bus avallon
					read 		<= 1'b1;
					byte_enable <= 4'hF;
                    // Le signal "acknoledge" est arrive, la lecture est terminee, on latch la donnee provenant du bus avallon pour la transmettre au bus SPI. 
                    if (ack_synchro) begin                      
                        reg_fstate [6:0]		<= 7'd4;
						read_data_to_spi[31:0] 	<= read_data_from_avallon_synchro[31:0];
					end
                    else begin
                        reg_fstate [6:0]	<= 7'd2;
						read_data_to_spi 	<= read_data_to_spi;
					end
                end
                7'd4: begin
                    // La lecture est terminee, les registres "read" et "byte_enable" sont remis a zero. On commence la transmission des donnees par le bus SPI. On attend le 64ieme bit pour passer a l'etat suivant.
					read 		<= 1'b0;            
					byte_enable <= 4'h0;
                    if (bit_cnt_synchro==7'h40)
                        reg_fstate [6:0] 	<= 7'd64;
                    else
                        reg_fstate [6:0] 	<= 7'd4;
                end
                7'd8: begin
                    // Debut de la reception de la donnee a ecrire en provenance du bus SPI. On attend le 64ieme bit pour passer a l'etat suivant : l'ecriture dans la memoire via le bus avallon.
                    if (bit_cnt_synchro==7'h40)
                        reg_fstate [6:0] 	<= 7'd16;
                    else
                        reg_fstate [6:0] 	<= 7'd8;
                end
                7'd16: begin
                    // Fin de la reception de la donnee, les registres "write" et "byte_enable" sont actif pour commencer l'operation d'ecriture.
                    // On inverse les octets de la donnee recue via le SPI
					write 					<= 1'b1;
					byte_enable 			<= 4'hF;
					write_data_to_avallon 	<= {data_from_spi_synchro[7:0], data_from_spi_synchro[15:8], data_from_spi_synchro[23:16], data_from_spi_synchro[31:24]};
                    if (ack_synchro)
                        reg_fstate [6:0] 	<= 7'd32;
                    else
                        reg_fstate [6:0] 	<= 7'd16;
                end
				7'd32: begin
                    // Le signal "csn" indique la fin de la trame, on retourne a l'etat IDLE
                    // Si l'on souhaite ecrire plusieurs donnees, on retourne a l'etat d'attente de la reception de la donnee SPI
					write 					<= 1'b0;
					byte_enable 			<= 4'h0;
					
					if (csn)
						reg_fstate [6:0] 	<= 7'd0;
					else if (bit_cnt_synchro==7'h20) begin
						reg_fstate [6:0] 	<= 7'd8;
						address 			<= address + 32'h1;
					end
					else
						reg_fstate [6:0] 	<= 7'd32;
				end
				7'd64: begin
                    // Comme pour l'etat precedent, le signal "csn" indique la fin de la trame, on retourne a l'etat IDLE
                    // Si l'on souhaite lire plusieurs donnees, on retourne a l'etat de demande de lecture au bus avallon
					if (csn)
						reg_fstate [6:0] 	<= 7'd0;
					else if (bit_cnt_synchro==7'h20) begin
						reg_fstate [6:0] 	<= 7'd2;
						address 			<= address + 32'h1;
					end
					else
						reg_fstate [6:0] 	<= 7'd64;
				end
                default: begin
					reg_fstate [6:0] 		<= 7'd0;
                end
            endcase
        end
    end
endmodule
